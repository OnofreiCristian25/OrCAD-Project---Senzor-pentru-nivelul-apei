** Profile: "SCHEMATIC1-simulare_oglinda"  [ c:\users\tedy_\desktop\pcad\proiect_oglinda-pspicefiles\schematic1\simulare_oglinda.sim ] 

** Creating circuit file "simulare_oglinda.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../mydiode.lib" 
* From [PSPICE NETLIST] section of C:\Users\Tedy_\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\22.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1000ns 0 
.STEP LIN PARAM r 28k 13k 100 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
